package dut_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "sequence_item.svh"

`include "reset_dut.svh"

`include "write_data.svh"
`include "read_data.svh"
`include "write_read.svh"
`include "wr_bulk.svh"
`include "write_err.svh"
`include "read_err.svh"


`include "driver.svh"

`include "result_monitor.svh"

`include "command_monitor.svh"


`include "agent.svh"

`include "scoreboard.svh"

`include "coverage.svh"

`include "env.svh"

`include "full_test.svh"


endpackage :dut_pkg
